module segLED (
	input [30:0] a,
	input [3:0] selin,
	output [7:0] out,
	output [3:0] sel
	);
	
	assign out = (a == 4'b0000) ? 8'b1111_1100:
					 (a == 4'b0001) ? 8'b0110_0000:
					 (a == 4'b0010) ? 8'b1101_1010:
					 (a == 4'b0011) ? 8'b1111_0010:
					 (a == 4'b0100) ? 8'b0110_0110:
					 (a == 4'b0101) ? 8'b1011_0110:
					 (a == 4'b0110) ? 8'b1011_1110:
					 (a == 4'b0111) ? 8'b1110_0000:
					 (a == 4'b1000) ? 8'b1111_1110:
					 (a == 4'b1001) ? 8'b1111_0110:
					 (a == 4'b1010) ? 8'b1110_1110:
				    (a == 4'b1011) ? 8'b0011_1110:
					 (a == 4'b1100) ? 8'b0001_1010:
					 (a == 4'b1101) ? 8'b0111_1010:
					 (a == 4'b1110) ? 8'b1001_1110:
					 8'b1000_1110;
	assign sel = selin;
endmodule