module shifter (
		input signed [15:0] A,
		input [3:0] opcode,
		input [3:0] d,
		output [15:0] Out,
		output [3:0] Outcond
		);
		wire [15:0] C;
		wire [15:0] D;
		wire [31:0] E;
		wire [3:0] cond;
		wire [0:0] cond1;
		assign D[15:0] = (opcode == 4'b1000) ? A << d:
							  (opcode == 4'b1001) ? C[15:0]:
							  (opcode == 4'b1010) ? A >> d:
							  A >>> d;
		assign E = A << d;
		assign C = (d == 4'b0000) ? E[15:0]:
					  (d == 4'b0001) ? {E[15:1],E[16]}:
					  (d == 4'b0010) ? {E[15:2],E[17:16]}:
					  (d == 4'b0011) ? {E[15:3],E[18:16]}:
					  (d == 4'b0100) ? {E[15:4],E[19:16]}:
					  (d == 4'b0101) ? {E[15:5],E[20:16]}:
					  (d == 4'b0110) ? {E[15:6],E[21:16]}:
					  (d == 4'b0111) ? {E[15:7],E[22:16]}:
					  (d == 4'b1000) ? {E[15:8],E[23:16]}:
					  (d == 4'b1001) ? {E[15:9],E[24:16]}:
					  (d == 4'b1010) ? {E[15:10],E[25:16]}:
					  (d == 4'b1011) ? {E[15:11],E[26:16]}:
					  (d == 4'b1100) ? {E[15:12],E[27:16]}:
					  (d == 4'b1101) ? {E[15:13],E[28:16]}:
					  (d == 4'b1110) ? {E[15:14],E[29:16]}:
					  {E[15],E[30:16]};
		assign cond1 = (d == 4'b0001) ? A[0]:
						   (d == 4'b0010) ? A[1]:
						   (d == 4'b0011) ? A[2]:
						   (d == 4'b0100) ? A[3]:
						   (d == 4'b0101) ? A[4]:
						   (d == 4'b0110) ? A[5]:
						   (d == 4'b0111) ? A[6]:
						   (d == 4'b1000) ? A[7]:
						   (d == 4'b1001) ? A[8]:
						   (d == 4'b1010) ? A[9]:
						   (d == 4'b1011) ? A[10]:
						   (d == 4'b1100) ? A[11]:
						   (d == 4'b1101) ? A[12]:
						   (d == 4'b1110) ? A[13]:
					      A[14];
		assign cond[0] = 1'b0;
		assign cond[1] = (d==0||opcode ==4'd9) ? 1'b0:
							  (opcode == 4'd8) ? E[16]:
							  cond1;
		assign cond[2] = (D[15:0]==16'b0) ? 1'b1:
							   1'b0;
		assign cond[3] = D[15];
		assign Out = D;
		assign Outcond = cond;
endmodule